package u8 is
  type unsigned8 is array (7 downto 0) of bit;
  type unsigned9 is array (8 downto 0) of bit;
end;
